`ifndef TRANSACTION
`define TRANSACTION

class transaction;
   bit reset;
  rand bit j;
  rand bit k;
  bit q;
  
endclass
`endif
